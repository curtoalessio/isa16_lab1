library verilog;
use verilog.vl_types.all;
entity tb_iir_adv is
end tb_iir_adv;
